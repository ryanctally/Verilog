module main;
  initial 
    begin
      $display("Learning Verilog is easy with referencedesigner.com tutorial");
      $finish ;
    end
endmodule
